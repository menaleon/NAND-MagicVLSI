magic
tech scmos
timestamp 1667975345
<< nwell >>
rect -13 2 26 22
<< polysilicon >>
rect -4 20 2 25
rect 11 20 17 25
rect -4 -7 2 3
rect 11 -7 17 3
rect -4 -29 2 -24
rect 11 -29 17 -24
<< ndiffusion >>
rect -12 -10 -4 -7
rect -12 -15 -11 -10
rect -6 -15 -4 -10
rect -12 -24 -4 -15
rect 2 -24 11 -7
rect 17 -10 25 -7
rect 17 -15 19 -10
rect 24 -15 25 -10
rect 17 -24 25 -15
<< pdiffusion >>
rect -12 10 -4 20
rect -12 5 -11 10
rect -6 5 -4 10
rect -12 3 -4 5
rect 2 10 11 20
rect 2 5 4 10
rect 9 5 11 10
rect 2 3 11 5
rect 17 10 25 20
rect 17 5 19 10
rect 24 5 25 10
rect 17 3 25 5
<< metal1 >>
rect -11 32 0 37
rect 5 32 24 37
rect -11 10 -6 32
rect 19 10 24 32
rect 4 -1 9 5
rect 4 -4 24 -1
rect 19 -10 24 -4
rect -11 -34 -6 -15
rect -11 -39 0 -34
rect 5 -39 13 -34
<< ntransistor >>
rect -4 -24 2 -7
rect 11 -24 17 -7
<< ptransistor >>
rect -4 3 2 20
rect 11 3 17 20
<< ndcontact >>
rect -11 -15 -6 -10
rect 19 -15 24 -10
<< pdcontact >>
rect -11 5 -6 10
rect 4 5 9 10
rect 19 5 24 10
<< nsubstratencontact >>
rect 0 32 5 37
rect 0 -39 5 -34
<< labels >>
rlabel polysilicon 1 -1 1 -1 1 a
rlabel polysilicon 12 -6 12 -6 1 b
rlabel metal1 7 -2 7 -2 1 out
rlabel metal1 9 34 9 34 5 vdd
rlabel metal1 8 -36 8 -36 1 gnd
<< end >>
