magic
tech scmos
timestamp 1667967760
<< nwell >>
rect -15 0 19 19
<< polysilicon >>
rect -4 18 -2 21
rect 7 18 9 21
rect -4 -9 -2 1
rect 7 -9 9 1
rect -4 -24 -2 -19
rect 7 -24 9 -19
<< ndiffusion >>
rect -14 -12 -4 -9
rect -14 -17 -12 -12
rect -7 -17 -4 -12
rect -14 -19 -4 -17
rect -2 -19 7 -9
rect 9 -12 18 -9
rect 9 -17 12 -12
rect 17 -17 18 -12
rect 9 -19 18 -17
<< pdiffusion >>
rect -14 12 -4 18
rect -14 7 -12 12
rect -7 7 -4 12
rect -14 1 -4 7
rect -2 12 7 18
rect -2 7 0 12
rect 5 7 7 12
rect -2 1 7 7
rect 9 12 18 18
rect 9 7 12 12
rect 17 7 18 12
rect 9 1 18 7
<< metal1 >>
rect -12 25 -4 30
rect 1 25 17 30
rect -12 12 -7 25
rect 12 12 17 25
rect 0 -3 5 7
rect 0 -6 17 -3
rect 12 -12 17 -6
rect -12 -28 -7 -17
rect -12 -32 -2 -28
rect 3 -32 9 -28
<< ntransistor >>
rect -4 -19 -2 -9
rect 7 -19 9 -9
<< ptransistor >>
rect -4 1 -2 18
rect 7 1 9 18
<< ndcontact >>
rect -12 -17 -7 -12
rect 12 -17 17 -12
<< pdcontact >>
rect -12 7 -7 12
rect 0 7 5 12
rect 12 7 17 12
<< nsubstratencontact >>
rect -4 25 1 30
rect -2 -32 3 -28
<< labels >>
rlabel polysilicon -3 -8 -3 -8 1 a
rlabel metal1 7 27 7 27 5 vdd
rlabel polysilicon 8 -7 8 -7 1 b
rlabel metal1 2 -3 2 -3 1 out
rlabel metal1 6 -30 6 -30 1 gnd
<< end >>
