* SPICE3 file created from nand_normal.ext - technology: scmos

.option scale=1u

M1000 vdd b out w_n13_2# pfet w=17 l=6
+  ad=272 pd=100 as=153 ps=52
M1001 out b a_2_n24# Gnd nfet w=17 l=6
+  ad=136 pd=50 as=153 ps=52
M1002 out a vdd w_n13_2# pfet w=17 l=6
+  ad=0 pd=0 as=0 ps=0
M1003 a_2_n24# a gnd Gnd nfet w=17 l=6
+  ad=0 pd=0 as=161 ps=70
C0 b w_n13_2# 2.14fF
C1 a w_n13_2# 2.14fF
C2 gnd 0 6.82fF **FLOATING
C3 out 0 3.38fF **FLOATING
C4 b 0 8.62fF **FLOATING
C5 a 0 8.62fF **FLOATING
C6 vdd 0 11.75fF **FLOATING
