* SPICE3 file created from nand_normal.ext - technology: scmos

.option scale=1u

.include ./ami05.txt
Vpower Vdd GND 5
Vin a gnd pulse(0,5,10n,1n,1n,10n,20n)
Vin2 b gnd pulse(0,5,10n,1n,10n,20n,20n)

M1000 vdd b out w_n10_2# pfet w=17 l=2
+  ad=306 pd=104 as=153 ps=52
M1001 out a vdd w_n10_2# pfet w=17 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out b a_2_n24# Gnd nfet w=17 l=2
+  ad=153 pd=52 as=153 ps=52
M1003 a_2_n24# a gnd Gnd nfet w=17 l=2
+  ad=0 pd=0 as=178 ps=72
C0 gnd 0 5.88fF 
C1 out 0 3.38fF 
C2 b 0 4.69fF 
C3 a 0 4.69fF 
C4 vdd 0 9.87fF 

.control 
run
set color0=white
set color1=black
set color2=blue
set color3=red
set xbrushwidth=5
plot a b out
.endc