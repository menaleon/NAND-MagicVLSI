magic
tech scmos
timestamp 1667964514
<< nwell >>
rect -10 2 23 14
<< polysilicon >>
rect 0 13 2 16
rect 11 13 13 16
rect 0 -7 2 3
rect 11 -7 13 3
rect 0 -22 2 -17
rect 11 -22 13 -17
<< ndiffusion >>
rect -9 -10 0 -7
rect -9 -15 -7 -10
rect -2 -15 0 -10
rect -9 -17 0 -15
rect 2 -17 11 -7
rect 13 -10 22 -7
rect 13 -15 15 -10
rect 20 -15 22 -10
rect 13 -17 22 -15
<< pdiffusion >>
rect -9 10 0 13
rect -9 5 -7 10
rect -2 5 0 10
rect -9 3 0 5
rect 2 10 11 13
rect 2 5 4 10
rect 9 5 11 10
rect 2 3 11 5
rect 13 10 22 13
rect 13 5 15 10
rect 20 5 22 10
rect 13 3 22 5
<< metal1 >>
rect -7 20 1 25
rect 6 20 20 25
rect -7 10 -2 20
rect 15 10 20 20
rect 4 -1 9 5
rect 4 -4 20 -1
rect 15 -10 20 -4
rect -7 -26 -2 -15
rect -7 -30 1 -26
rect 6 -30 13 -26
<< ntransistor >>
rect 0 -17 2 -7
rect 11 -17 13 -7
<< ptransistor >>
rect 0 3 2 13
rect 11 3 13 13
<< ndcontact >>
rect -7 -15 -2 -10
rect 15 -15 20 -10
<< pdcontact >>
rect -7 5 -2 10
rect 4 5 9 10
rect 15 5 20 10
<< nsubstratencontact >>
rect 1 20 6 25
rect 1 -30 6 -26
<< labels >>
rlabel metal1 9 -28 9 -28 1 gnd
rlabel polysilicon 1 -1 1 -1 1 a
rlabel polysilicon 12 -6 12 -6 1 b
rlabel metal1 11 23 11 23 5 vdd
rlabel metal1 7 -2 7 -2 1 out
<< end >>
