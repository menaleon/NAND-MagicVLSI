* SPICE3 file created from nand_normal.ext - technology: scmos

.option scale=1u

M1000 vdd b out w_n10_2# pfet w=17 l=2
+  ad=306 pd=104 as=153 ps=52
M1001 out a vdd w_n10_2# pfet w=17 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out b a_2_n24# Gnd nfet w=17 l=2
+  ad=153 pd=52 as=153 ps=52
M1003 a_2_n24# a gnd Gnd nfet w=17 l=2
+  ad=0 pd=0 as=178 ps=72
C0 gnd 0 5.88fF **FLOATING
C1 out 0 3.38fF **FLOATING
C2 b 0 4.69fF **FLOATING
C3 a 0 4.69fF **FLOATING
C4 vdd 0 9.87fF **FLOATING
