* SPICE3 file created from nand_normal.ext - technology: scmos

.option scale=1u

.include ./ami05.txt
Vpower Vdd GND 5
Vin a gnd pulse(0,5,10n,1n,1n,10n,20n)
Vin2 b gnd pulse(0,5,10n,1n,10n,20n,20n)

M1000 a_2_n17# a gnd Gnd nfet w=10 l=2
+  ad=90 pd=38 as=110 ps=56
M1001 vdd b out w_n12_2# pfet w=10 l=6
+  ad=160 pd=72 as=70 ps=34
M1002 out b a_2_n17# Gnd nfet w=10 l=2
+  ad=90 pd=38 as=0 ps=0
M1003 out a vdd w_n12_2# pfet w=10 l=6
+  ad=0 pd=0 as=0 ps=0
C0 gnd 0 4.93fF 
C1 out 0 3.38fF 
C2 b 0 5.56fF 
C3 a 0 5.56fF 
C4 vdd 0 8.93fF 

.control 
run
set color0=white
set color1=black
set color2=blue
set color3=red
set xbrushwidth=5
plot a b out
.endc
.tran 0.01 40n
.end