magic
tech scmos
timestamp 1667972284
<< nwell >>
rect -11 6 22 18
<< polysilicon >>
rect -1 17 1 20
rect 10 17 12 20
rect -1 -3 1 7
rect 10 -3 12 7
rect -1 -25 1 -20
rect 10 -25 12 -20
<< ndiffusion >>
rect -10 -11 -1 -3
rect -10 -16 -8 -11
rect -3 -16 -1 -11
rect -10 -20 -1 -16
rect 1 -20 10 -3
rect 12 -11 21 -3
rect 12 -16 14 -11
rect 19 -16 21 -11
rect 12 -20 21 -16
<< pdiffusion >>
rect -10 14 -1 17
rect -10 9 -8 14
rect -3 9 -1 14
rect -10 7 -1 9
rect 1 14 10 17
rect 1 9 3 14
rect 8 9 10 14
rect 1 7 10 9
rect 12 14 21 17
rect 12 9 14 14
rect 19 9 21 14
rect 12 7 21 9
<< metal1 >>
rect -8 24 0 29
rect 5 24 19 29
rect -8 14 -3 24
rect 14 14 19 24
rect 3 3 8 9
rect 3 0 19 3
rect 14 -11 19 0
rect -8 -29 -3 -16
rect -8 -33 0 -29
rect 5 -33 12 -29
<< ntransistor >>
rect -1 -20 1 -3
rect 10 -20 12 -3
<< ptransistor >>
rect -1 7 1 17
rect 10 7 12 17
<< ndcontact >>
rect -8 -16 -3 -11
rect 14 -16 19 -11
<< pdcontact >>
rect -8 9 -3 14
rect 3 9 8 14
rect 14 9 19 14
<< nsubstratencontact >>
rect 0 24 5 29
rect 0 -33 5 -29
<< labels >>
rlabel metal1 10 27 10 27 5 vdd
rlabel metal1 5 3 5 3 1 out
rlabel polysilicon 0 0 0 0 1 a
rlabel polysilicon 11 -1 11 -1 1 b
rlabel metal1 8 -31 8 -31 1 gnd
<< end >>
