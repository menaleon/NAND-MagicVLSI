magic
tech scmos
timestamp 1667973694
<< nwell >>
rect -12 2 25 14
<< polysilicon >>
rect -3 13 3 16
rect 10 13 16 16
rect -3 1 3 3
rect 10 1 16 3
rect 0 -7 2 1
rect 11 -7 13 1
rect 0 -22 2 -17
rect 11 -22 13 -17
<< ndiffusion >>
rect -9 -10 0 -7
rect -9 -15 -7 -10
rect -2 -15 0 -10
rect -9 -17 0 -15
rect 2 -17 11 -7
rect 13 -10 22 -7
rect 13 -15 15 -10
rect 20 -15 22 -10
rect 13 -17 22 -15
<< pdiffusion >>
rect -11 10 -3 13
rect -11 5 -9 10
rect -4 5 -3 10
rect -11 3 -3 5
rect 3 10 10 13
rect 3 5 4 10
rect 9 5 10 10
rect 3 3 10 5
rect 16 10 24 13
rect 16 5 17 10
rect 22 5 24 10
rect 16 3 24 5
<< metal1 >>
rect -9 20 1 25
rect 6 20 22 25
rect -9 10 -4 20
rect 17 10 22 20
rect 4 -1 9 5
rect 4 -4 20 -1
rect 15 -10 20 -4
rect -7 -26 -2 -15
rect -7 -30 1 -26
rect 6 -30 13 -26
<< ntransistor >>
rect 0 -17 2 -7
rect 11 -17 13 -7
<< ptransistor >>
rect -3 3 3 13
rect 10 3 16 13
<< ndcontact >>
rect -7 -15 -2 -10
rect 15 -15 20 -10
<< pdcontact >>
rect -9 5 -4 10
rect 4 5 9 10
rect 17 5 22 10
<< nsubstratencontact >>
rect 1 20 6 25
rect 1 -30 6 -26
<< labels >>
rlabel metal1 9 -28 9 -28 1 gnd
rlabel polysilicon 1 -1 1 -1 1 a
rlabel polysilicon 12 -6 12 -6 1 b
rlabel metal1 11 23 11 23 5 vdd
rlabel metal1 7 -2 7 -2 1 out
<< end >>
