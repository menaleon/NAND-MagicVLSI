* SPICE3 file created from nand_normal.ext - technology: scmos

.option scale=1u

M1000 vdd b out w_n10_2# pfet w=10 l=2
+  ad=180 pd=76 as=90 ps=38
M1001 out a vdd w_n10_2# pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out b a_3_n17# Gnd nfet w=10 l=6
+  ad=90 pd=38 as=70 ps=34
M1003 a_3_n17# a gnd Gnd nfet w=10 l=6
+  ad=0 pd=0 as=110 ps=56
C0 gnd 0 5.50fF **FLOATING
C1 out 0 3.81fF **FLOATING
C2 b 0 6.82fF **FLOATING
C3 a 0 6.82fF **FLOATING
C4 vdd 0 7.99fF **FLOATING
