* SPICE3 file created from nand_aumentoWn.ext - technology: scmos

.option scale=1u

M1000 a_1_n20# a gnd Gnd nfet w=17 l=2
+  ad=153 pd=52 as=173 ps=70
M1001 out a vdd w_n11_6# pfet w=10 l=2
+  ad=90 pd=38 as=180 ps=76
M1002 out b a_1_n20# Gnd nfet w=17 l=2
+  ad=153 pd=52 as=0 ps=0
M1003 vdd b out w_n11_6# pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd 0 4.93fF **FLOATING
C1 out 0 3.38fF **FLOATING
C2 b 0 4.45fF **FLOATING
C3 a 0 4.45fF **FLOATING
C4 vdd 0 7.99fF **FLOATING
