magic
tech scmos
timestamp 1667974879
<< nwell >>
rect -10 2 23 22
<< polysilicon >>
rect 0 20 2 25
rect 11 20 13 25
rect 0 -7 2 3
rect 11 -7 13 3
rect 0 -29 2 -24
rect 11 -29 13 -24
<< ndiffusion >>
rect -9 -10 0 -7
rect -9 -15 -7 -10
rect -2 -15 0 -10
rect -9 -24 0 -15
rect 2 -24 11 -7
rect 13 -10 22 -7
rect 13 -15 15 -10
rect 20 -15 22 -10
rect 13 -24 22 -15
<< pdiffusion >>
rect -9 10 0 20
rect -9 5 -7 10
rect -2 5 0 10
rect -9 3 0 5
rect 2 10 11 20
rect 2 5 4 10
rect 9 5 11 10
rect 2 3 11 5
rect 13 10 22 20
rect 13 5 15 10
rect 20 5 22 10
rect 13 3 22 5
<< metal1 >>
rect -7 32 0 37
rect 5 32 20 37
rect -7 10 -2 32
rect 15 10 20 32
rect 4 -1 9 5
rect 4 -4 20 -1
rect 15 -10 20 -4
rect -7 -34 -2 -15
rect -7 -39 0 -34
rect 5 -39 13 -34
<< ntransistor >>
rect 0 -24 2 -7
rect 11 -24 13 -7
<< ptransistor >>
rect 0 3 2 20
rect 11 3 13 20
<< ndcontact >>
rect -7 -15 -2 -10
rect 15 -15 20 -10
<< pdcontact >>
rect -7 5 -2 10
rect 4 5 9 10
rect 15 5 20 10
<< nsubstratencontact >>
rect 0 32 5 37
rect 0 -39 5 -34
<< labels >>
rlabel polysilicon 1 -1 1 -1 1 a
rlabel polysilicon 12 -6 12 -6 1 b
rlabel metal1 7 -2 7 -2 1 out
rlabel metal1 9 34 9 34 5 vdd
rlabel metal1 8 -36 8 -36 1 gnd
<< end >>
