magic
tech scmos
timestamp 1667976125
<< nwell >>
rect -13 2 26 13
<< polysilicon >>
rect -4 13 2 18
rect 11 13 17 18
rect -4 -7 2 3
rect 11 -7 17 3
rect -4 -20 2 -17
rect 11 -20 17 -17
<< ndiffusion >>
rect -12 -9 -4 -7
rect -12 -14 -11 -9
rect -6 -14 -4 -9
rect -12 -17 -4 -14
rect 2 -17 11 -7
rect 17 -9 25 -7
rect 17 -14 19 -9
rect 24 -14 25 -9
rect 17 -17 25 -14
<< pdiffusion >>
rect -12 10 -4 13
rect -12 5 -11 10
rect -6 5 -4 10
rect -12 3 -4 5
rect 2 10 11 13
rect 2 5 4 10
rect 9 5 11 10
rect 2 3 11 5
rect 17 10 25 13
rect 17 5 19 10
rect 24 5 25 10
rect 17 3 25 5
<< metal1 >>
rect -11 23 -3 28
rect 2 23 24 28
rect -11 10 -6 23
rect 19 10 24 23
rect 4 -1 9 5
rect 4 -4 24 -1
rect 19 -9 24 -4
rect -11 -29 -6 -14
rect -11 -34 -4 -29
rect 1 -34 17 -29
<< ntransistor >>
rect -4 -17 2 -7
rect 11 -17 17 -7
<< ptransistor >>
rect -4 3 2 13
rect 11 3 17 13
<< ndcontact >>
rect -11 -14 -6 -9
rect 19 -14 24 -9
<< pdcontact >>
rect -11 5 -6 10
rect 4 5 9 10
rect 19 5 24 10
<< nsubstratencontact >>
rect -3 23 2 28
rect -4 -34 1 -29
<< labels >>
rlabel polysilicon 1 -1 1 -1 1 a
rlabel polysilicon 12 -6 12 -6 1 b
rlabel metal1 7 -2 7 -2 1 out
rlabel metal1 12 26 12 26 5 vdd
rlabel metal1 7 -31 7 -31 1 gnd
<< end >>
