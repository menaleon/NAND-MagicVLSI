* SPICE3 file created from nand_normal.ext - technology: scmos

.option scale=1u

M1000 vdd b out w_n10_2# pfet w=10 l=2
+  ad=180 pd=76 as=90 ps=38
M1001 a_2_n17# a gnd Gnd nfet w=10 l=2
+  ad=90 pd=38 as=110 ps=56
M1002 out a vdd w_n10_2# pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out b a_2_n17# Gnd nfet w=10 l=2
+  ad=90 pd=38 as=0 ps=0
C0 gnd 0 4.93fF **FLOATING
C1 out 0 3.38fF **FLOATING
C2 b 0 4.45fF **FLOATING
C3 a 0 4.45fF **FLOATING
C4 vdd 0 7.99fF **FLOATING
